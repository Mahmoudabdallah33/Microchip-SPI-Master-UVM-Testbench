package spi_master_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "spi_master_seq_item.sv"
`include "spi_master_sqr.sv"
`include "spi_master_agt_config.sv"
`include "spi_master_env_config.sv"

`include "spi_master_seq.sv"
`include "spi_master_drv.sv"
`include "spi_master_mon.sv"

`include "spi_master_agt.sv"
`include "spi_master_cov.sv"
`include "spi_master_predictor.sv"
`include "spi_master_evaluator.sv"
`include "spi_master_scb.sv"
`include "spi_master_env.sv"
`include "spi_test.sv"



endpackage
