class spi_master_sqr extends uvm_sequencer #(spi_master_seq_item);
   `uvm_component_utils(spi_master_sqr)
  function new(string name = "spi_master_sqr",uvm_component parent);
   super.new(name,parent);
 
  endfunction 

  




endclass
